module main

pub fn optimize(node Node) Node {
	return node
}
