module ske

pub fn optimize(node Node) Node {
	return node
}
