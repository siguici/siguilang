module eval

import ske.ast
import ske.checker { is_bool, is_float, is_int }

pub struct Var {
pub mut:
	type    Type
	value   Value
	mutable bool
}

pub struct Eval {
mut:
	vars map[string]Var
	ctx  Context
}

pub fn Eval.new() Eval {
	return Eval{}
}

pub fn new_eval() Eval {
	return Eval.new()
}

pub fn eval(program ast.Program) ! {
	mut ev := new_eval()
	ev.eval(program)!
}

pub fn (mut this Eval) init_var(type string, name string, value Value) ! {
	var_type := Type.from(type)
	is_valid := if value !is Nil && var_type is BuiltinType {
		(var_type.is(.bool) && value.is_bool())
			|| (var_type.is(.int) && value.is_int())
			|| (var_type.is(.float) && value.is_float())
			|| (var_type.is(.string) && value.is_string())
	} else {
		true
	}
	if !is_valid {
		return error('Invalid type for variable ${name} (got ${value.type_name()} expected ${type})')
	} else {
		this.vars[name] = Var{
			type:    Type.from(type)
			value:   value
			mutable: name.starts_with('\$')
		}
	}
}

pub fn (mut this Eval) set_var(name string, value Value) ! {
	if var_def := this.vars[name] {
		if !var_def.mutable {
			return error('Cannot modify read-only variable ${name}')
		}
		this.vars[name].value = value
	} else {
		return error('Undefined variable ${name}')
	}
}

pub fn (this Eval) get_var(name string) !Value {
	return if var_def := this.vars[name] {
		var_def.value
	} else {
		error('Undefined variable ${name}')
	}
}

pub fn (mut this Eval) eval(p ast.Program) ! {
	for node in p.nodes {
		this.eval_node(node)!
	}
}

pub fn (mut this Eval) eval_node(n ast.Node) ! {
	match n {
		ast.Block {
			this.eval_block(n)!
		}
		ast.Stmt {
			this.eval_stmt(n)!
		}
		ast.EmptyNode {
			this.eval_empty(n)
		}
	}
}
